library ieee;
use ieee.std_logic_1164.all;

entity constants is
	port(s: IN std_logic;
		a : IN std_logic_vector(7 downto 0);
		oprnd: OUT std_logic_vector(7 downto 0));
end constants;

architecture beh of constants is
begin
	process(s,a)
	begin
		if(s='0')then
			oprnd<="ZZZZZZZZ";
		elsif(s='1')then
			oprnd<=a;
		end if;
	end process;
end beh;